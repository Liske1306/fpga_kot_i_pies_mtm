module char_rom_16x16
    (
        input  logic       clk,
        input  logic [7:0] char_xy,            // {x[3:0], y[3:0]}
        output logic [6:0]  char_code // pixels of the character line
    );

    logic [6:0] text[0:15][0:15] = '{{7'h64, 7'h62, 7'h72, 7'h62, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h01},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h61, 7'h62, 7'h72, 7'h61, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h62},
    {7'h63, 7'h62, 7'h72, 7'h62, 7'h6B, 7'h61, 7'h64, 7'h61, 7'h62, 7'h72, 7'h61, 7'h61, 7'h61, 7'h61, 7'h61, 7'h68} 
    };

    always_ff @(posedge clk) begin
        char_code <= text[char_xy[3:0]][char_xy[7:4]];
    end

endmodule